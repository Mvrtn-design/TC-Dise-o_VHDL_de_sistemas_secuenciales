library ieee;  
use ieee.std_logic_1164.all;

entity practica_2 is
port (clk, rst, x: in std_logic;
z: out std_logic);
end practica_2;